module ball (
	input wire clk,
	input wire reset,
	input wire [19:0] paddle_state,
	output reg [19:0] ball_pos,
	output reg [1:0] score_state
);
	

endmodule
