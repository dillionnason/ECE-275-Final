module score (
	input wire reset,
	input wire [1:0] score_state,
	output reg [5:0] current_score,
	output reg game_over
);

endmodule
